LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY int7seg IS
	PORT (
		d : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		dOut : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END int7seg;

ARCHITECTURE logicFunction OF int7seg IS

	SIGNAL Ndout : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

	dOut <= "11000000" WHEN d = "0000" ELSE
		"11111001" WHEN d = "0001" ELSE
		"10100100" WHEN d = "0010" ELSE
		"10110000" WHEN d = "0011" ELSE
		"10011001" WHEN d = "0100" ELSE
		"10010010" WHEN d = "0101" ELSE
		"10000010" WHEN d = "0110" ELSE
		"11111000" WHEN d = "0111" ELSE
		"10000000" WHEN d = "1000" ELSE
		"10011000" WHEN d = "1001" ELSE
		"10001000" WHEN d = "1010" ELSE
		"10000011" WHEN d = "1011" ELSE
		"11000110" WHEN d = "1100" ELSE
		"10100001" WHEN d = "1101" ELSE
		"10000110" WHEN d = "1110" ELSE
		"10001110";

END LogicFunction;